`ifndef DEFS_SVH
`define DEFS_SVH

`define XLEN 32
`define NUM_REGS 32

`define BYTE_WIDTH 8
`define INST_WIDTH 32

`endif